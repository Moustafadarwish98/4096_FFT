// ============================================================================
// Purpose:
//   Performs Bit-Reversal Reordering for a streaming FFT.
//
// Description:
//   In a Decimation-in-Frequency (DIF) FFT, outputs naturally emerge in
//   bit-reversed order. This module buffers the entire frame and reads it
//   back using bit-reversed addressing so that samples exit in natural order.
//
// Operation:
//   1. Incoming samples are written sequentially into memory (wraddr).
//   2. Read address (rdaddr) is generated by reversing wraddr bits.
//   3. MSB is inverted to ensure correct double-buffering behavior.
//   4. After one full frame is written, outputs become valid.
// ============================================================================

`default_nettype none

module bitreverse #(
    // ------------------------------------------------------------------------
    // Configuration Parameters
    // ------------------------------------------------------------------------
    parameter LGSIZE = 5,   // log2(FFT size / samples per frame)
    parameter WIDTH  = 24   // Bit width of each complex sample
)(
    // ------------------------------------------------------------------------
    // Ports
    // ------------------------------------------------------------------------
    input  wire                 i_clk,
    input  wire                 i_reset,
    input  wire                 i_clk_enable,

    input  wire [(2*WIDTH-1):0] i_in,    // Complex input sample
    output reg  [(2*WIDTH-1):0] o_out,   // Bit-reversed output
    output reg                  o_sync   // Output frame sync
);

  // ========================================================================
  // 1. ADDRESS GENERATION
  // ========================================================================
  //
  // wraddr:
  //   Sequential write pointer.
  //   Width = LGSIZE+1 to support frame toggling (MSB = bank select).
  //
  // rdaddr:
  //   Bit-reversed version of wraddr.
  //   Used to read memory in natural FFT order.

  reg  [(LGSIZE):0] wraddr;
  wire [(LGSIZE):0] rdaddr;

  // ========================================================================
  // 2. MEMORY BUFFER
  // ========================================================================
  //
  // brmem:
  //   Dual-frame buffer (size = 2^(LGSIZE+1)).
  //   Stores an entire FFT frame before valid readout begins.
  //
  // Why double size?
  //   MSB of wraddr acts as a "ping-pong" bank selector so that
  //   reading and writing can occur without collision.

  reg [(2*WIDTH-1):0] brmem [0:((1<<(LGSIZE))-1)];

  // ========================================================================
  // 3. BIT-REVERSED READ ADDRESS
  // ========================================================================
  //
  // rdaddr[k] = reversed(wraddr[k])
  //
  // Example (LGSIZE=4):
  //   wraddr = b3 b2 b1 b0
  //   rdaddr = b0 b1 b2 b3
  //
  // This mapping restores natural FFT bin order.

  genvar k;
  generate
    for (k = 0; k < LGSIZE; k = k + 1)
    begin : GEN_BIT_REVERSE
      assign rdaddr[k] = wraddr[LGSIZE-1-k];
    end
  endgenerate

  // MSB inversion:
  //   Toggles between memory banks.
  //   Ensures correct pipeline scheduling.

  assign rdaddr[LGSIZE] = !wraddr[LGSIZE];

  // ========================================================================
  // 4. RESET TRACKING (VALIDITY CONTROL)
  // ========================================================================
  //
  // in_reset:
  //   Remains high until one full frame has been written.
  //
  // Why needed?
  //   Prevents asserting o_sync while memory still contains invalid data.

  reg in_reset;

  always @(posedge i_clk)
    if (i_reset)
      in_reset <= 1'b1;
    else if ((i_clk_enable) && (&wraddr[(LGSIZE-1):0]))
      // All lower bits = 1 → End of frame reached
      in_reset <= 1'b0;

  // ========================================================================
  // 5. WRITE LOGIC (INPUT BUFFERING)
  // ========================================================================
  //
  // Stores incoming samples sequentially.
  //
  // wraddr increments every enabled clock.
  // Memory depth supports full-frame buffering.

  always @(posedge i_clk)
    if (i_reset)
      wraddr <= 0;
    else if (i_clk_enable)
    begin
      brmem[wraddr] <= i_in;  // Store sample
      wraddr <= wraddr + 1;   // Advance pointer
    end

  // ========================================================================
  // 6. READ LOGIC (BIT-REVERSED OUTPUT)
  // ========================================================================
  //
  // Reads memory using rdaddr.
  //
  // Note:
  //   No explicit reset condition needed.
  //   Invalid outputs during reset are ignored via o_sync gating.

  always @(posedge i_clk)
    if (i_clk_enable)
      o_out <= brmem[rdaddr];

  // ========================================================================
  // 7. OUTPUT SYNC GENERATION
  // ========================================================================
  //
  // o_sync asserted at start of each valid output frame.
  //
  // Condition:
  //   wraddr lower bits == 0 → First sample of frame
  //   AND not in_reset → Memory now contains valid FFT data

  always @(posedge i_clk)
    if (i_reset)
      o_sync <= 1'b0;
    else if ((i_clk_enable) && (!in_reset))
      o_sync <= (wraddr[(LGSIZE-1):0] == 0);

endmodule
