`include "register_interface/typedef.svh"
`include "register_interface/assign.svh"

module butterfly_top #(
    parameter int unsigned AXI_ADDR_WIDTH = 32,
    localparam int unsigned AXI_DATA_WIDTH = 32,
    parameter int unsigned AXI_ID_WIDTH = -1,
    parameter int unsigned AXI_USER_WIDTH = -1
)(
    input  logic          clk_i,
    input  logic          rst_ni,
    input  logic          test_mode_i,
    AXI_BUS.Slave         axi_slave
);

    // Import the types autogenerated by reggen
    import butterfly_reg_pkg::butterfly_reg2hw_t;
    import butterfly_reg_pkg::butterfly_hw2reg_t;

    // Declare the internal Register Bus interface
    REG_BUS #(
        .ADDR_WIDTH(32),
        .DATA_WIDTH(32)
    ) axi_to_regfile();
    // =========================================================================
    // STEP 3.5: Declare Register-to-Hardware and Hardware-to-Register Wires
    // =========================================================================
    // These structs represent the physical wires connecting the autogenerated
    // register file to your custom butterfly IP. 
    // They are typed using the imports we declared at the top of the module.
    
    // Carries operands and control signals from software to hardware
    butterfly_reg2hw_t reg_file_to_ip;  
    
    // Carries results and status flags from hardware back to software
    butterfly_hw2reg_t ip_to_reg_file;  


    // =========================================================================
    // STEP 3.6: Instantiate the AXI-to-Register Protocol Converter
    // =========================================================================
    // The PULP SoC uses the AXI protocol, but our autogenerated register file 
    // uses a simpler Generic Register Protocol. 
    // This module acts as the bridge, converting AXI transactions on `axi_slave` 
    // into register read/write transactions on `axi_to_regfile`.
    
    axi_to_reg_intf #(
        .ADDR_WIDTH (AXI_ADDR_WIDTH),
        .DATA_WIDTH (AXI_DATA_WIDTH),
        .ID_WIDTH   (AXI_ID_WIDTH),
        .USER_WIDTH (AXI_USER_WIDTH),
        .DECOUPLE_W (0)
    ) i_axi2reg (
        .clk_i      (clk_i),
        .rst_ni     (rst_ni),
        .testmode_i (test_mode_i),
        .in         (axi_slave),      // The AXI port exposed to the SoC crossbar
        .reg_o      (axi_to_regfile)  // The internal REG_BUS interface
    );


    // =========================================================================
    // STEP 3.7: Convert the REG_BUS Interface to Reggen Structs
    // =========================================================================
    // The autogenerated register file doesn't use SystemVerilog interfaces.
    // It expects flat structs for requests and responses. These macros handle
    // the conversion smoothly without introducing logic delays.

    // 1. Define the basic types matching AXI widths
    typedef logic [AXI_ADDR_WIDTH-1:0]   addr_t;
    typedef logic [AXI_DATA_WIDTH-1:0]   data_t;
    typedef logic [AXI_DATA_WIDTH/8-1:0] strb_t;

// 2. Use PULP macros to create the request/response struct types
    `REG_BUS_TYPEDEF_REQ(reg_req_t, addr_t, data_t, strb_t)
    `REG_BUS_TYPEDEF_RSP(reg_rsp_t, data_t)

    // 3. Declare the actual struct wires
    reg_req_t to_reg_file_req;   
    reg_rsp_t from_reg_file_rsp; 

    // 4. Map the signals between the REG_BUS interface and the structs
    `REG_BUS_ASSIGN_TO_REQ(to_reg_file_req, axi_to_regfile)
    `REG_BUS_ASSIGN_FROM_RSP(axi_to_regfile, from_reg_file_rsp)
    // =========================================================================
    // STEP 3.8: Instantiate the Autogenerated Register File
    // =========================================================================
    // This is the module generated by the reggen tool. It takes the converted 
    // struct requests (from Step 3.7) and exposes the physical hardware wires.
    
    butterfly_reg_top #(
        .reg_req_t(reg_req_t),
        .reg_rsp_t(reg_rsp_t)
    ) i_regfile (
        .clk_i      (clk_i),
        .rst_ni     (rst_ni),
        .devmode_i  (1'b1), // Tied to 1 for standalone IPs as per PULP convention
        
        // From AXI-to-register protocol converter
        .reg_req_i  (to_reg_file_req),
        .reg_rsp_o  (from_reg_file_rsp),
        
        // Connections to the Butterfly IP
        .reg2hw     (reg_file_to_ip),
        .hw2reg     (ip_to_reg_file)
    );

    // =========================================================================
    // STEP 3.9: Instantiate and Wire the Butterfly Accelerator
    // =========================================================================
    
    // Intermediate wires for outputs to safely map to multireg structs
    logic [37:0] butterfly_o_left;
    logic [37:0] butterfly_o_right;
    logic        butterfly_o_aux;

    // Instance of the actual Hardware Accelerator
    butterfly #(
        .IWIDTH(19),
        .CWIDTH(23),
        .OWIDTH(19),
        .SHIFT(0),
        .CKPCE(1)
    ) i_butterfly (
        .i_clk        (clk_i),
        .i_reset      (~rst_ni),
        
        // --- Control Signals ---
        // .q holds the stable value, .qe pulses high for 1 cycle on write
        .i_clk_enable (reg_file_to_ip.ctrl.enable.q),
        .i_aux        (reg_file_to_ip.ctrl.trigger.q & reg_file_to_ip.ctrl.trigger.qe),
        
        // --- Input Operands (Unpacking from multireg arrays) ---
        // Coef is 46 bits: [1] holds upper 14 bits, [0] holds lower 32 bits
        .i_coef       ({reg_file_to_ip.coef[1].q[13:0], reg_file_to_ip.coef[0].q}),
        
        // Left/Right inputs are 38 bits: [1] holds upper 6 bits, [0] holds lower 32 bits
        .i_left       ({reg_file_to_ip.op_left[1].q[5:0], reg_file_to_ip.op_left[0].q}),
        .i_right      ({reg_file_to_ip.op_right[1].q[5:0], reg_file_to_ip.op_right[0].q}),
        
        // --- Outputs ---
        .o_left       (butterfly_o_left),
        .o_right      (butterfly_o_right),
        .o_aux        (butterfly_o_aux)
    );

    // --- Output Mapping (Packing into multireg arrays) ---
    // When o_aux pulses high, the hardware writes the results back to the registers
    
// Status DONE bit
    assign ip_to_reg_file.status.d  = 1'b1;             
    assign ip_to_reg_file.status.de = butterfly_o_aux;

    // Result Left
    assign ip_to_reg_file.result_left[0].d  = butterfly_o_left[31:0];
    assign ip_to_reg_file.result_left[1].d  = {26'b0, butterfly_o_left[37:32]};
    assign ip_to_reg_file.result_left[0].de = butterfly_o_aux; 
    assign ip_to_reg_file.result_left[1].de = butterfly_o_aux;

    // Result Right
    assign ip_to_reg_file.result_right[0].d  = butterfly_o_right[31:0];
    assign ip_to_reg_file.result_right[1].d  = {26'b0, butterfly_o_right[37:32]};
    assign ip_to_reg_file.result_right[0].de = butterfly_o_aux;
    assign ip_to_reg_file.result_right[1].de = butterfly_o_aux;
    
    // Hardware Diagnostic Prints
    always @(posedge clk_i) begin
        if (reg_file_to_ip.ctrl.trigger.q & reg_file_to_ip.ctrl.trigger.qe)
            $display("[HW DEBUG] CYCLE %0t: AXI Trigger received! i_aux is HIGH", $time);
            
        if (butterfly_o_aux)
            $display("[HW DEBUG] CYCLE %0t: Pipeline Finished! o_aux is HIGH", $time);
    end

endmodule
